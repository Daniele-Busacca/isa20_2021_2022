library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IMEM_ABS is
    generic( m : positive := 30;       -- ADD parallelism
             n : positive := 32);     -- DOUT parallelism
    port (
        ADD : in std_logic_vector( m-1 downto 0 );
        -------------------------------------------
        DOUT : out std_logic_vector( n-1 downto 0 )
    );
end IMEM_ABS;

architecture beh of IMEM_ABS is

    type MEM_Array is array ( 0 to 25 ) of std_logic_vector( n-1 downto 0 );

    signal MEM : MEM_Array := ( "00000000011100000000100000010011",
                                "00001111110000010000001000010111",
                                "11111111110000100000001000010011",
                                "00001111110000010000001010010111",
                                "00000001000000101000001010010011",
                                "01000000000000000000011010110111",
                                "11111111111101101000011010010011",
                                "00000010000010000000100001100011",
                                "00000000000000100010010000000011",
                                "01000000000001000001010100100000",
                                "00000000000000000000000000000000",
                                "00000000000000000000000000000000",
                                "00000000000000000000000000000000",
                                "00000000010000100000001000010011",
                                "11111111111110000000100000010011",
                                "00000000110101010010010110110011",
                                "11111100000001011000111011100011",
                                "00000000000001010000011010110011",
                                "11111101010111111111000011101111",
                                "00000000110100101010000000100011",
                                "00000000000000000000000011101111",
                                "00000000000000000000000000010011",
                                "00000000000000000000000000000000",
                                "00000000000000000000000000000000",
                                "00000000000000000000000000000000",
                                "00000000000000000000000000000000"
                                );

                                
    begin

        MEM_Process : process( ADD )

        begin

            DOUT <= MEM(to_integer(unsigned(ADD)));
        
        end process;


end architecture;
