library ieee;
use ieee.std_logic_1164.all;

entity Dec5to32 is
    port (
        A : in std_logic_vector( 4 downto 0 );
        ---------------------------------------
        Y : out std_logic_vector( 31 downto 0 )
    );
end Dec5to32;

architecture beh of Dec5to32 is

    begin

        Y <= "00000000000000000000000000000001" when A = "00000" else
             "00000000000000000000000000000010" when A = "00001" else
             "00000000000000000000000000000100" when A = "00010" else
             "00000000000000000000000000001000" when A = "00011" else
             "00000000000000000000000000010000" when A = "00100" else
             "00000000000000000000000000100000" when A = "00101" else
             "00000000000000000000000001000000" when A = "00110" else
             "00000000000000000000000010000000" when A = "00111" else
             "00000000000000000000000100000000" when A = "01000" else
             "00000000000000000000001000000000" when A = "01001" else
             "00000000000000000000010000000000" when A = "01010" else
             "00000000000000000000100000000000" when A = "01011" else
             "00000000000000000001000000000000" when A = "01100" else
             "00000000000000000010000000000000" when A = "01101" else
             "00000000000000000100000000000000" when A = "01110" else
             "00000000000000001000000000000000" when A = "01111" else
             "00000000000000010000000000000000" when A = "10000" else
             "00000000000000100000000000000000" when A = "10001" else
             "00000000000001000000000000000000" when A = "10010" else
             "00000000000010000000000000000000" when A = "10011" else
             "00000000000100000000000000000000" when A = "10100" else
             "00000000001000000000000000000000" when A = "10101" else
             "00000000010000000000000000000000" when A = "10110" else
             "00000000100000000000000000000000" when A = "10111" else
             "00000001000000000000000000000000" when A = "11000" else
             "00000010000000000000000000000000" when A = "11001" else
             "00000100000000000000000000000000" when A = "11010" else
             "00001000000000000000000000000000" when A = "11011" else
             "00010000000000000000000000000000" when A = "11100" else
             "00100000000000000000000000000000" when A = "11101" else
             "01000000000000000000000000000000" when A = "11110" else
             "10000000000000000000000000000000";

end architecture;